// Copyright 2022 Intel Corporation
// SPDX-License-Identifier: MIT

`ifndef dma_vh

    `define dma_vh
    
    `define DMA_DO_SINGLE_BURST_PARTIAL_WRITES 1

`endif
