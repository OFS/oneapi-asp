// Copyright 2020 Intel Corporation.
//
// THIS SOFTWARE MAY CONTAIN PREPRODUCTION CODE AND IS PROVIDED BY THE
// COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED
// WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
// MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR
// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,
// WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE
// OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE,
// EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//

`include "ofs_plat_if.vh"
`include "opencl_bsp.vh"


module afu
import dc_bsp_pkg::*;
  #(
    parameter NUM_LOCAL_MEM_BANKS = 0,
    parameter NUM_ETH = 0
   )
  (
    // Host memory (Avalon)
    ofs_plat_avalon_mem_rdwr_if.to_sink host_mem_if,

    // FPGA MMIO master (Avalon)
    ofs_plat_avalon_mem_if.to_source mmio64_if,

    // Local memory interface.
    ofs_plat_avalon_mem_if.to_slave local_mem[NUM_LOCAL_MEM_BANKS],
    
    `ifdef INCLUDE_UDP_OFFLOAD_ENGINE
        // Ethernet
        ofs_fim_hssi_ss_tx_axis_if.client eth_tx_axis ,
        ofs_fim_hssi_ss_rx_axis_if.client eth_rx_axis ,
        ofs_fim_hssi_fc_if.client     eth_fc ,
    `endif

    // clocks and reset
    input logic pClk,                      //Primary interface clock
    input logic pClk_reset,                // ACTIVE HIGH Soft Reset
    input logic uClk_usr,                  // User clock domain. Refer to clock programming guide
    input logic uClk_usr_reset,
    input logic uClk_usrDiv2,              // User clock domain. Half the programmed frequency
    input logic uClk_usrDiv2_reset
);

import dma_pkg::*;

logic reset, clk;
assign reset = pClk_reset;
assign clk   = pClk;

//local wires to connect between bsp_logic and kernel_wrapper - kernel control and memory-interface
opencl_kernel_control_intf opencl_kernel_control();
kernel_mem_intf kernel_mem[BSP_NUM_LOCAL_MEM_BANKS]();

`ifdef USE_MPF_VTP
    // The width of the Avalon-MM user field is narrower on the AFU side
    // of VTP, since VTP uses a bit to flag VTP page table traffic.
    // Drop the high bit of the user field on the AFU side.
    localparam AFU_AVMM_USER_WIDTH = host_mem_if.USER_WIDTH_ - 1;
    
    // Virtual address interface for use by the DMA path.
    ofs_plat_avalon_mem_rdwr_if
    #(
        `OFS_PLAT_AVALON_MEM_RDWR_IF_REPLICATE_PARAMS_EXCEPT_TAGS(host_mem_if),
        .USER_WIDTH(AFU_AVMM_USER_WIDTH),
        .LOG_CLASS(ofs_plat_log_pkg::HOST_CHAN)
    ) host_mem_va_if();
    
    assign host_mem_va_if.clk = host_mem_if.clk;
    assign host_mem_va_if.reset_n = host_mem_if.reset_n;
    assign host_mem_va_if.instance_number = host_mem_if.instance_number;
    
    // mmio64-if for the BSP
    ofs_plat_avalon_mem_if
    #(
        `OFS_PLAT_AVALON_MEM_IF_REPLICATE_PARAMS(mmio64_if)
    ) mmio64_if_shim();
    
    assign mmio64_if_shim.clk = mmio64_if.clk;
    assign mmio64_if_shim.reset_n = mmio64_if.reset_n;
    assign mmio64_if_shim.instance_number = mmio64_if.instance_number;
    
    mem_if_vtp mem_if_vtp_inst (
        .host_mem_if,
        .host_mem_va_if,
        .mmio64_if,
        .mmio64_if_shim
    );
`endif

`ifdef INCLUDE_UDP_OFFLOAD_ENGINE
//UDP/HSSI offload engine
    shim_avst_if udp_avst_from_kernel();
    shim_avst_if udp_avst_to_kernel();
    ofs_plat_avalon_mem_if #(
        `OFS_PLAT_AVALON_MEM_IF_REPLICATE_PARAMS(mmio64_if)
    ) uoe_csr_avmm();
    assign uoe_csr_avmm.clk     = clk;
    assign uoe_csr_avmm.reset_n = ~reset;
    
    udp_offload_engine udp_offload_engine
    (
        //MAC interfaces
        .eth_rx_axis,
        .eth_tx_axis,
        .eth_fc,
    
        // kernel clock and reset
        .kernel_clk(uClk_usrDiv2),
        .kernel_resetn(opencl_kernel_control.kernel_reset_n),
    
        // from kernel
        .udp_avst_from_kernel,
        
        // to kernel
        .udp_avst_to_kernel,
    
        // CSR
        .uoe_csr_avmm
    );
`endif

//BSP/shim logic

bsp_logic bsp_logic_inst (
    .clk                    ( pClk ),
    .reset,
    .kernel_clk             ( uClk_usrDiv2 ),
    .kernel_clk_reset       ( uClk_usrDiv2_reset ),
    `ifdef USE_MPF_VTP
        .host_mem_if        ( host_mem_va_if ),
        .mmio64_if          ( mmio64_if_shim ),
    `else
        .host_mem_if        ( host_mem_if ),
        .mmio64_if          ( mmio64_if ),
    `endif
    `ifdef INCLUDE_UDP_OFFLOAD_ENGINE
        .uoe_csr_avmm,
    `endif
    .local_mem,
    
    .opencl_kernel_control,
    .kernel_mem
);

kernel_wrapper kernel_wrapper_inst (
    .clk        (uClk_usrDiv2),
    .clk2x      (uClk_usr),
    .reset_n    (!uClk_usrDiv2_reset),
    .opencl_kernel_control,
    .kernel_mem
`ifdef INCLUDE_USM_SUPPORT
    , .kernel_svm           ( host_mem_pa_if_kernel )
`endif
`ifdef INCLUDE_UDP_OFFLOAD_ENGINE
    ,.udp_avst_from_kernel,
    .udp_avst_to_kernel
`endif
);

endmodule : afu
